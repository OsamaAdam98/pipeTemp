`include "pipeTemp.v"

module pipeTempTest;

    pipeTemp PipeTemp(8'd100);

endmodule