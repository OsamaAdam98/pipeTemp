`include "pipeTemp.v"

module pipeTempTest;

    pipeTemp PipeTemp(8'd200);

endmodule